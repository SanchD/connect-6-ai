module controller(
	input clk,
	input reset,
	input data_in,
	output data_out
	);

endmodule